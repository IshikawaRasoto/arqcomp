library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity calculadora is
    port(
        entrada: in std_logic,
        saida: out std_logic
    );
end entity;
    